library verilog;
use verilog.vl_types.all;
entity test_cache is
end test_cache;
